module	lcd_run (
					iCLK,	
start,enable,
					LCD_DATA,LCD_RW,LCD_EN,LCD_RS, select_lcd);
input [3:0] select_lcd;
input			iCLK;
input start,enable;
output	[7:0]	LCD_DATA;
output			LCD_RW,LCD_EN,LCD_RS;
reg	[5:0]	LUT_INDEX;
reg	[8:0]	LUT_DATA;
reg	[5:0]	mLCD_ST;
reg	[17:0]	mDLY;
reg			mLCD_Start;
reg	[7:0]	mLCD_DATA;
reg			mLCD_RS;
wire		mLCD_Done;
wire clk_out;
parameter	LCD_INTIAL	=	0;
parameter	LCD_LINE1	=	5;
parameter	LCD_CH_LINE	=	LCD_LINE1+16;
parameter	LCD_LINE2	=	LCD_LINE1+16+1;
parameter	LUT_SIZE	=	LCD_LINE1+32+1;
div_to_1 clock_out(.CLOCK_50(iCLK),.clk_out(clk_out));
always@(posedge iCLK /*or negedge clk_out*/)
begin
	if(!1)
	begin
		LUT_INDEX	<=	0;
		mLCD_ST		<=	0;
		mDLY			<=	0;
		mLCD_Start	<=	0;
		mLCD_DATA	<=	0;
		mLCD_RS		<=	0;
	end
	else
	begin
		if(LUT_INDEX<LUT_SIZE)
		begin
			case(mLCD_ST)
			0:	begin
					mLCD_DATA	<=	LUT_DATA[7:0];
					mLCD_RS		<=	LUT_DATA[8];
					mLCD_Start	<=	1;
					mLCD_ST		<=	1;
				end
			1:	begin
					if(mLCD_Done)
					begin
						mLCD_Start	<=	0;
						mLCD_ST		<=	2;					
					end
				end
			2:	begin
					if(mDLY<18'h3FFFE)
					mDLY	<=	mDLY+1;
					else
					begin
						mDLY	<=	0;
						mLCD_ST	<=	3;
						
					end
				end
			3:	begin
					LUT_INDEX	<=	LUT_INDEX+1;
					mLCD_ST	<=	0;
				end
			endcase
		end
		else LUT_INDEX<=LCD_LINE1;
	end
end

always
begin
case(select_lcd)
	4'b0001: 
	begin
	case(LUT_INDEX)
	//	Initial
	LCD_INTIAL+0:	LUT_DATA	<=	9'h038;
	LCD_INTIAL+1:	LUT_DATA	<=	9'h00C;
	LCD_INTIAL+2:	LUT_DATA	<=	9'h001;
	LCD_INTIAL+3:	LUT_DATA	<=	9'h006;
	LCD_INTIAL+4:	LUT_DATA	<=	9'h080;
	//	Line 1
	LCD_LINE1+0:	LUT_DATA	<=	9'h120;	//_!!ALERT-ON!!__
	LCD_LINE1+1:	LUT_DATA	<=	9'h120;
	LCD_LINE1+2:	LUT_DATA	<=	9'h121; //!
	LCD_LINE1+3:	LUT_DATA	<=	9'h121; //!
	LCD_LINE1+4:	LUT_DATA	<=	9'h141; //A
	LCD_LINE1+5:	LUT_DATA	<=	9'h14C; //L
	LCD_LINE1+6:	LUT_DATA	<=	9'h145; //E
	LCD_LINE1+7:	LUT_DATA	<=	9'h152; //R
	LCD_LINE1+8:	LUT_DATA	<=	9'h154; //T
	LCD_LINE1+9:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE1+10:	LUT_DATA	<=	9'h14F; //O
	LCD_LINE1+11:	LUT_DATA	<=	9'h14E; //N
	LCD_LINE1+12:	LUT_DATA	<=	9'h121; //!
	LCD_LINE1+13:	LUT_DATA	<=	9'h121; //!
	LCD_LINE1+14:	LUT_DATA	<=	9'h120;
	LCD_LINE1+15:	LUT_DATA	<=	9'h120;
	//	Change Line
	LCD_CH_LINE:	LUT_DATA	<=	9'h0C0;
	//	Line 2
	LCD_LINE2+0:	LUT_DATA	<=	9'h120;	//_!!ALERT-ON!!__
	LCD_LINE2+1:	LUT_DATA	<=	9'h120;
	LCD_LINE2+2:	LUT_DATA	<=	9'h121; //!
	LCD_LINE2+3:	LUT_DATA	<=	9'h121; //!
	LCD_LINE2+4:	LUT_DATA	<=	9'h141; //A
	LCD_LINE2+5:	LUT_DATA	<=	9'h14C; //L
	LCD_LINE2+6:	LUT_DATA	<=	9'h145; //E
	LCD_LINE2+7:	LUT_DATA	<=	9'h152; //R
	LCD_LINE2+8:	LUT_DATA	<=	9'h154; //T
	LCD_LINE2+9:	LUT_DATA	<= 9'h15F; //- 
	LCD_LINE2+10:	LUT_DATA	<=	9'h14F; //O
	LCD_LINE2+11:	LUT_DATA	<=	9'h14E; //N
	LCD_LINE2+12:	LUT_DATA	<=	9'h121; //!
	LCD_LINE2+13:	LUT_DATA	<=	9'h121; //!
	LCD_LINE2+14:	LUT_DATA	<=	9'h120;
	LCD_LINE2+15:	LUT_DATA	<=	9'h120;
	default:		LUT_DATA	<=	9'h120;
	endcase
	end
	4'b0010: 
	begin
	case(LUT_INDEX)
	//	Initial
	LCD_INTIAL+0:	LUT_DATA	<=	9'h038;
	LCD_INTIAL+1:	LUT_DATA	<=	9'h00C;
	LCD_INTIAL+2:	LUT_DATA	<=	9'h001;
	LCD_INTIAL+3:	LUT_DATA	<=	9'h006;
	LCD_INTIAL+4:	LUT_DATA	<=	9'h080;
	//	Line 1
	LCD_LINE1+0:	LUT_DATA	<=	9'h120;	//_!!ALERT-OFF!!_
	LCD_LINE1+1:	LUT_DATA	<=	9'h120;
	LCD_LINE1+2:	LUT_DATA	<=	9'h121; //!
	LCD_LINE1+3:	LUT_DATA	<=	9'h121; //!
	LCD_LINE1+4:	LUT_DATA	<=	9'h141; //A
	LCD_LINE1+5:	LUT_DATA	<=	9'h14C; //L
	LCD_LINE1+6:	LUT_DATA	<=	9'h145; //E
	LCD_LINE1+7:	LUT_DATA	<=	9'h152; //R
	LCD_LINE1+8:	LUT_DATA	<=	9'h154; //T
	LCD_LINE1+9:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE1+10:	LUT_DATA	<=	9'h14F; //O
	LCD_LINE1+11:	LUT_DATA	<=	9'h146; //F
	LCD_LINE1+12:	LUT_DATA	<=	9'h146; //F
	LCD_LINE1+13:	LUT_DATA	<=	9'h121; //!
	LCD_LINE1+14:	LUT_DATA	<=	9'h121; //!
	LCD_LINE1+15:	LUT_DATA	<=	9'h120;
	//	Change Line
	LCD_CH_LINE:	LUT_DATA	<=	9'h0C0;
	//	Line 2
	LCD_LINE2+0:	LUT_DATA	<=	9'h120;	//_!!ALERT-OFF!!_
	LCD_LINE2+1:	LUT_DATA	<=	9'h120;
	LCD_LINE2+2:	LUT_DATA	<=	9'h121; //!
	LCD_LINE2+3:	LUT_DATA	<=	9'h121; //!
	LCD_LINE2+4:	LUT_DATA	<=	9'h141; //A
	LCD_LINE2+5:	LUT_DATA	<=	9'h14C; //L
	LCD_LINE2+6:	LUT_DATA	<=	9'h145; //E
	LCD_LINE2+7:	LUT_DATA	<=	9'h152; //R
	LCD_LINE2+8:	LUT_DATA	<=	9'h154; //T
	LCD_LINE2+9:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE2+10:	LUT_DATA	<=	9'h14F; //O
	LCD_LINE2+11:	LUT_DATA	<=	9'h146; //F
	LCD_LINE2+12:	LUT_DATA	<=	9'h146; //F
	LCD_LINE2+13:	LUT_DATA	<=	9'h121; //!
	LCD_LINE2+14:	LUT_DATA	<=	9'h121; //!
	LCD_LINE2+15:	LUT_DATA	<=	9'h120;
	default:		LUT_DATA	<=	9'h120;
	endcase
	end
	4'b0011: 
	begin
	case(LUT_INDEX)
	//	Initial
	LCD_INTIAL+0:	LUT_DATA	<=	9'h038;
	LCD_INTIAL+1:	LUT_DATA	<=	9'h00C;
	LCD_INTIAL+2:	LUT_DATA	<=	9'h001;
	LCD_INTIAL+3:	LUT_DATA	<=	9'h006;
	LCD_INTIAL+4:	LUT_DATA	<=	9'h080;
	//	Line 1
	LCD_LINE1+0:	LUT_DATA	<=	9'h120;	//_<FINDINGCAR>_
	LCD_LINE1+1:	LUT_DATA	<=	9'h120;
	LCD_LINE1+2:	LUT_DATA	<=	9'h13C; //<
	LCD_LINE1+3:	LUT_DATA	<=	9'h146; //F
	LCD_LINE1+4:	LUT_DATA	<=	9'h149; //I
	LCD_LINE1+5:	LUT_DATA	<=	9'h14E; //N
	LCD_LINE1+6:	LUT_DATA	<=	9'h144; //D
	LCD_LINE1+7:	LUT_DATA	<=	9'h149; //I
	LCD_LINE1+8:	LUT_DATA	<=	9'h14E; //N
	LCD_LINE1+9:	LUT_DATA	<=	9'h147; //G
	LCD_LINE1+10:	LUT_DATA	<=	9'h143; //C
	LCD_LINE1+11:	LUT_DATA	<=	9'h141; //A
	LCD_LINE1+12:	LUT_DATA	<=	9'h152; //R
	LCD_LINE1+13:	LUT_DATA	<=	9'h13E; //>
	LCD_LINE1+14:	LUT_DATA	<=	9'h120; 
	LCD_LINE1+15:	LUT_DATA	<=	9'h120;
	//	Change Line
	LCD_CH_LINE:	LUT_DATA	<=	9'h0C0;
	//	Line 2
	LCD_LINE2+0:	LUT_DATA	<=	9'h120;	//_<FINDINGCAR>_
	LCD_LINE2+1:	LUT_DATA	<=	9'h120;
	LCD_LINE2+2:	LUT_DATA	<=	9'h13C; //<
	LCD_LINE2+3:	LUT_DATA	<=	9'h146; //F
	LCD_LINE2+4:	LUT_DATA	<=	9'h149; //I
	LCD_LINE2+5:	LUT_DATA	<=	9'h14E; //N
	LCD_LINE2+6:	LUT_DATA	<=	9'h144; //D
	LCD_LINE2+7:	LUT_DATA	<=	9'h149; //I
	LCD_LINE2+8:	LUT_DATA	<=	9'h14E; //N
	LCD_LINE2+9:	LUT_DATA	<=	9'h147; //G
	LCD_LINE2+10:	LUT_DATA	<=	9'h143; //C
	LCD_LINE2+11:	LUT_DATA	<=	9'h141; //A
	LCD_LINE2+12:	LUT_DATA	<=	9'h152; //R
	LCD_LINE2+13:	LUT_DATA	<=	9'h13E; //>
	LCD_LINE2+14:	LUT_DATA	<=	9'h120; 
	LCD_LINE2+15:	LUT_DATA	<=	9'h120;
	default:		LUT_DATA	<=	9'h120;
	endcase
	end
	4'b0100: 
	begin
	case(LUT_INDEX)
	//	Initial
	LCD_INTIAL+0:	LUT_DATA	<=	9'h038;
	LCD_INTIAL+1:	LUT_DATA	<=	9'h00C;
	LCD_INTIAL+2:	LUT_DATA	<=	9'h001;
	LCD_INTIAL+3:	LUT_DATA	<=	9'h006;
	LCD_INTIAL+4:	LUT_DATA	<=	9'h080;
	//	Line 1
	LCD_LINE1+0:	LUT_DATA	<=	9'h120;	//_<VERIFYPASS>_
	LCD_LINE1+1:	LUT_DATA	<=	9'h120;
	LCD_LINE1+2:	LUT_DATA	<=	9'h13C; //<
	LCD_LINE1+3:	LUT_DATA	<=	9'h156; //V
	LCD_LINE1+4:	LUT_DATA	<=	9'h145; //E
	LCD_LINE1+5:	LUT_DATA	<=	9'h152; //R
	LCD_LINE1+6:	LUT_DATA	<=	9'h149; //I
	LCD_LINE1+7:	LUT_DATA	<=	9'h146; //F
	LCD_LINE1+8:	LUT_DATA	<=	9'h159; //Y
	LCD_LINE1+9:	LUT_DATA	<=	9'h150; //P
	LCD_LINE1+10:	LUT_DATA	<=	9'h141; //A
	LCD_LINE1+11:	LUT_DATA	<=	9'h153; //S
	LCD_LINE1+12:	LUT_DATA	<=	9'h153; //S
	LCD_LINE1+13:	LUT_DATA	<=	9'h13E; //>
	LCD_LINE1+14:	LUT_DATA	<=	9'h120; 
	LCD_LINE1+15:	LUT_DATA	<=	9'h120;
	//	Change Line
	LCD_CH_LINE:	LUT_DATA	<=	9'h0C0;
	//	Line 2
	LCD_LINE2+0:	LUT_DATA	<=	9'h120;	//_<PASS-WRONG>__
	LCD_LINE2+1:	LUT_DATA	<=	9'h120;
	LCD_LINE2+2:	LUT_DATA	<=	9'h13C; //<
	LCD_LINE2+3:	LUT_DATA	<=	9'h150; //P
	LCD_LINE2+4:	LUT_DATA	<=	9'h141; //A
	LCD_LINE2+5:	LUT_DATA	<=	9'h153; //S
	LCD_LINE2+6:	LUT_DATA	<=	9'h153; //S
	LCD_LINE2+7:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE2+8:	LUT_DATA	<=	9'h157; //W
	LCD_LINE2+9:	LUT_DATA	<=	9'h152; //R
	LCD_LINE2+10:	LUT_DATA	<=	9'h14F; //O
	LCD_LINE2+11:	LUT_DATA	<=	9'h14E; //N
	LCD_LINE2+12:	LUT_DATA	<=	9'h147; //G
	LCD_LINE2+13:	LUT_DATA	<=	9'h13E; //>
	LCD_LINE2+14:	LUT_DATA	<=	9'h120; 
	LCD_LINE2+15:	LUT_DATA	<=	9'h120;
	default:		LUT_DATA	<=	9'h120;
	endcase
	end
	4'b0101: 
	begin
	case(LUT_INDEX)
	//	Initial
	LCD_INTIAL+0:	LUT_DATA	<=	9'h038;
	LCD_INTIAL+1:	LUT_DATA	<=	9'h00C;
	LCD_INTIAL+2:	LUT_DATA	<=	9'h001;
	LCD_INTIAL+3:	LUT_DATA	<=	9'h006;
	LCD_INTIAL+4:	LUT_DATA	<=	9'h080;
	//	Line 1
	LCD_LINE1+0:	LUT_DATA	<=	9'h120;	//_<VERIFYPASS>_
	LCD_LINE1+1:	LUT_DATA	<=	9'h120;
	LCD_LINE1+2:	LUT_DATA	<=	9'h13C; //<
	LCD_LINE1+3:	LUT_DATA	<=	9'h156; //V
	LCD_LINE1+4:	LUT_DATA	<=	9'h145; //E
	LCD_LINE1+5:	LUT_DATA	<=	9'h152; //R
	LCD_LINE1+6:	LUT_DATA	<=	9'h149; //I
	LCD_LINE1+7:	LUT_DATA	<=	9'h146; //F
	LCD_LINE1+8:	LUT_DATA	<=	9'h159; //Y
	LCD_LINE1+9:	LUT_DATA	<=	9'h150; //P
	LCD_LINE1+10:	LUT_DATA	<=	9'h141; //A
	LCD_LINE1+11:	LUT_DATA	<=	9'h153; //S
	LCD_LINE1+12:	LUT_DATA	<=	9'h153; //S
	LCD_LINE1+13:	LUT_DATA	<=	9'h13E; //>
	LCD_LINE1+14:	LUT_DATA	<=	9'h120; 
	LCD_LINE1+15:	LUT_DATA	<=	9'h120;
	//	Change Line
	LCD_CH_LINE:	LUT_DATA	<=	9'h0C0;
	//	Line 2
	LCD_LINE2+0:	LUT_DATA	<=	9'h120;	//_<PASS-RIGHT>__
	LCD_LINE2+1:	LUT_DATA	<=	9'h120;
	LCD_LINE2+2:	LUT_DATA	<=	9'h13C; //<
	LCD_LINE2+3:	LUT_DATA	<=	9'h150; //P
	LCD_LINE2+4:	LUT_DATA	<=	9'h141; //A
	LCD_LINE2+5:	LUT_DATA	<=	9'h153; //S
	LCD_LINE2+6:	LUT_DATA	<=	9'h153; //S
	LCD_LINE2+7:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE2+8:	LUT_DATA	<=	9'h152; //R
	LCD_LINE2+9:	LUT_DATA	<=	9'h149; //I
	LCD_LINE2+10:	LUT_DATA	<=	9'h147; //G
	LCD_LINE2+11:	LUT_DATA	<=	9'h148; //H
	LCD_LINE2+12:	LUT_DATA	<=	9'h154; //T
	LCD_LINE2+13:	LUT_DATA	<=	9'h13E; //>
	LCD_LINE2+14:	LUT_DATA	<=	9'h120; 
	LCD_LINE2+15:	LUT_DATA	<=	9'h120;
	default:		LUT_DATA	<=	9'h120;
	endcase
	end
	4'b0110: 
	begin
	case(LUT_INDEX)
	//	Initial
	LCD_INTIAL+0:	LUT_DATA	<=	9'h038;
	LCD_INTIAL+1:	LUT_DATA	<=	9'h00C;
	LCD_INTIAL+2:	LUT_DATA	<=	9'h001;
	LCD_INTIAL+3:	LUT_DATA	<=	9'h006;
	LCD_INTIAL+4:	LUT_DATA	<=	9'h080;
	//	Line 1
	LCD_LINE1+0:	LUT_DATA	<=	9'h120;	//_<VERIFYPASS>_
	LCD_LINE1+1:	LUT_DATA	<=	9'h120;
	LCD_LINE1+2:	LUT_DATA	<=	9'h13C; //<
	LCD_LINE1+3:	LUT_DATA	<=	9'h156; //V
	LCD_LINE1+4:	LUT_DATA	<=	9'h145; //E
	LCD_LINE1+5:	LUT_DATA	<=	9'h152; //R
	LCD_LINE1+6:	LUT_DATA	<=	9'h149; //I
	LCD_LINE1+7:	LUT_DATA	<=	9'h146; //F
	LCD_LINE1+8:	LUT_DATA	<=	9'h159; //Y
	LCD_LINE1+9:	LUT_DATA	<=	9'h150; //P
	LCD_LINE1+10:	LUT_DATA	<=	9'h141; //A
	LCD_LINE1+11:	LUT_DATA	<=	9'h153; //S
	LCD_LINE1+12:	LUT_DATA	<=	9'h153; //S
	LCD_LINE1+13:	LUT_DATA	<=	9'h13E; //>
	LCD_LINE1+14:	LUT_DATA	<=	9'h120; 
	LCD_LINE1+15:	LUT_DATA	<=	9'h120;
	//	Change Line
	LCD_CH_LINE:	LUT_DATA	<=	9'h0C0;
	//	Line 2
	LCD_LINE2+0:	LUT_DATA	<=	9'h120;	//_<VERIFYPASS>_
	LCD_LINE2+1:	LUT_DATA	<=	9'h120;
	LCD_LINE2+2:	LUT_DATA	<=	9'h13C; //<
	LCD_LINE2+3:	LUT_DATA	<=	9'h156; //V
	LCD_LINE2+4:	LUT_DATA	<=	9'h145; //E
	LCD_LINE2+5:	LUT_DATA	<=	9'h152; //R
	LCD_LINE2+6:	LUT_DATA	<=	9'h149; //I
	LCD_LINE2+7:	LUT_DATA	<=	9'h146; //F
	LCD_LINE2+8:	LUT_DATA	<=	9'h159; //Y
	LCD_LINE2+9:	LUT_DATA	<=	9'h150; //P
	LCD_LINE2+10:	LUT_DATA	<=	9'h141; //A
	LCD_LINE2+11:	LUT_DATA	<=	9'h153; //S
	LCD_LINE2+12:	LUT_DATA	<=	9'h153; //S
	LCD_LINE2+13:	LUT_DATA	<=	9'h13E; //>
	LCD_LINE2+14:	LUT_DATA	<=	9'h120; 
	LCD_LINE2+15:	LUT_DATA	<=	9'h120;
	default:		LUT_DATA	<=	9'h120;
	endcase
	end
	4'b0111: 
	begin
	case(LUT_INDEX)
	//	Initial
	LCD_INTIAL+0:	LUT_DATA	<=	9'h038;
	LCD_INTIAL+1:	LUT_DATA	<=	9'h00C;
	LCD_INTIAL+2:	LUT_DATA	<=	9'h001;
	LCD_INTIAL+3:	LUT_DATA	<=	9'h006;
	LCD_INTIAL+4:	LUT_DATA	<=	9'h080;
	//	Line 1
	LCD_LINE1+0:	LUT_DATA	<=	9'h120;	//_---START--->_
	LCD_LINE1+1:	LUT_DATA	<=	9'h120;
	LCD_LINE1+2:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE1+3:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE1+4:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE1+5:	LUT_DATA	<=	9'h153; //S
	LCD_LINE1+6:	LUT_DATA	<=	9'h154; //T
	LCD_LINE1+7:	LUT_DATA	<=	9'h141; //A
	LCD_LINE1+8:	LUT_DATA	<=	9'h152; //R
	LCD_LINE1+9:	LUT_DATA	<=	9'h154; //T
	LCD_LINE1+10:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE1+11:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE1+12:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE1+13:	LUT_DATA	<=	9'h13E; //>
	LCD_LINE1+14:	LUT_DATA	<=	9'h120; 
	LCD_LINE1+15:	LUT_DATA	<=	9'h120;
	//	Change Line
	LCD_CH_LINE:	LUT_DATA	<=	9'h0C0;
	//	Line 2
	LCD_LINE2+0:	LUT_DATA	<=	9'h120;	//_---START--->_
	LCD_LINE2+1:	LUT_DATA	<=	9'h120;
	LCD_LINE2+2:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE2+3:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE2+4:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE2+5:	LUT_DATA	<=	9'h153; //S
	LCD_LINE2+6:	LUT_DATA	<=	9'h154; //T
	LCD_LINE2+7:	LUT_DATA	<=	9'h141; //A
	LCD_LINE2+8:	LUT_DATA	<=	9'h152; //R
	LCD_LINE2+9:	LUT_DATA	<=	9'h154; //T
	LCD_LINE2+10:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE2+11:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE2+12:	LUT_DATA	<=	9'h15F; //-
	LCD_LINE2+13:	LUT_DATA	<=	9'h13E; //>
	LCD_LINE2+14:	LUT_DATA	<=	9'h120; 
	LCD_LINE2+15:	LUT_DATA	<=	9'h120;
	default:		LUT_DATA	<=	9'h120;
	endcase
	end
	4'b0000:
	begin
	case(LUT_INDEX)
	//	Initial
	LCD_INTIAL+0:	LUT_DATA	<=	9'h038;
	LCD_INTIAL+1:	LUT_DATA	<=	9'h00C;
	LCD_INTIAL+2:	LUT_DATA	<=	9'h001;
	LCD_INTIAL+3:	LUT_DATA	<=	9'h006;
	LCD_INTIAL+4:	LUT_DATA	<=	9'h080;
	//	Line 1
	/*LCD_LINE1+0:	LUT_DATA	<=	9'h120;	//_[]BLOCKCAR[]_
	LCD_LINE1+1:	LUT_DATA	<=	9'h120;
	LCD_LINE1+2:	LUT_DATA	<=	9'h15B; //[
	LCD_LINE1+3:	LUT_DATA	<=	9'h15D; //]
	LCD_LINE1+4:	LUT_DATA	<=	9'h142; //B
	LCD_LINE1+5:	LUT_DATA	<=	9'h14C; //L
	LCD_LINE1+6:	LUT_DATA	<=	9'h14F; //O
	LCD_LINE1+7:	LUT_DATA	<=	9'h143; //C
	LCD_LINE1+8:	LUT_DATA	<=	9'h14B; //K
	LCD_LINE1+9:	LUT_DATA	<=	9'h143; //C
	LCD_LINE1+10:	LUT_DATA	<=	9'h141; //A
	LCD_LINE1+11:	LUT_DATA	<=	9'h152; //R
	LCD_LINE1+12:	LUT_DATA	<=	9'h15B; //[
	LCD_LINE1+13:	LUT_DATA	<=	9'h15D; //]
	LCD_LINE1+14:	LUT_DATA	<=	9'h120; 
	LCD_LINE1+15:	LUT_DATA	<=	9'h120;*/
	
	LCD_LINE1+0:	LUT_DATA	<=	9'h120;	
	LCD_LINE1+1:	LUT_DATA	<=	9'h120;
	LCD_LINE1+2:	LUT_DATA	<=	9'h120;
	LCD_LINE1+3:	LUT_DATA	<=	9'h143; //C
	LCD_LINE1+4:	LUT_DATA	<= 9'h141; //A
	LCD_LINE1+5:	LUT_DATA	<=	9'h152; //R
	LCD_LINE1+6:	LUT_DATA	<=	9'h12D; //-
	LCD_LINE1+7:	LUT_DATA	<=	9'h153; //S
	LCD_LINE1+8:	LUT_DATA	<=	9'h154; //T
	LCD_LINE1+9:	LUT_DATA	<=	9'h141; //A
	LCD_LINE1+10:	LUT_DATA	<=	9'h154; //T
	LCD_LINE1+11:	LUT_DATA	<=	9'h145; //E
	LCD_LINE1+12:	LUT_DATA	<=	9'h13A; //:
	LCD_LINE1+13:	LUT_DATA	<=	9'h120;
	LCD_LINE1+14:	LUT_DATA	<=	9'h120; 
	LCD_LINE1+15:	LUT_DATA	<=	9'h120;
	//	Change Line
	LCD_CH_LINE:	LUT_DATA	<=	9'h0C0;
	//	Line 2
	LCD_LINE2+0:	LUT_DATA	<=	9'h120;	//_[]BLOCKCAR[]_
	LCD_LINE2+1:	LUT_DATA	<=	9'h120;
	LCD_LINE2+2:	LUT_DATA	<=	9'h15B; //[
	LCD_LINE2+3:	LUT_DATA	<=	9'h15D; //]
	LCD_LINE2+4:	LUT_DATA	<=	9'h142; //B
	LCD_LINE2+5:	LUT_DATA	<=	9'h14C; //L
	LCD_LINE2+6:	LUT_DATA	<=	9'h14F; //O
	LCD_LINE2+7:	LUT_DATA	<=	9'h143; //C
	LCD_LINE2+8:	LUT_DATA	<=	9'h14B; //K
	LCD_LINE2+9:	LUT_DATA	<=	9'h143; //C
	LCD_LINE2+10:	LUT_DATA	<=	9'h141; //A
	LCD_LINE2+11:	LUT_DATA	<=	9'h152; //R
	LCD_LINE2+12:	LUT_DATA	<=	9'h15B; //[
	LCD_LINE2+13:	LUT_DATA	<=	9'h15D; //]
	LCD_LINE2+14:	LUT_DATA	<=	9'h120; 
	LCD_LINE2+15:	LUT_DATA	<=	9'h120;
	default:		LUT_DATA	<=	9'h120;
	endcase
	end
endcase
end

LCD_Controller u0	(
							.iDATA(mLCD_DATA),
							.iRS(mLCD_RS),
							.iStart(mLCD_Start),
							.oDone(mLCD_Done),
							.iCLK(iCLK),
							.start(start),
							.LCD_DATA(LCD_DATA),
							.LCD_RW(LCD_RW),
							.LCD_EN(LCD_EN),
							.LCD_RS(LCD_RS)	);

endmodule

