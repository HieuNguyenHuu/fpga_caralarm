module car-test();





car (CLOCK_50 ,LCD_DATA, LCD_RW, LCD_RS, LCD_EN,IRDA_RXD,
SW,KEY,HEX0,HEX1,HEX2,HEX3,HEX4,HEX5,HEX6,HEX7,LEDR,LEDG);



















endmodule 


